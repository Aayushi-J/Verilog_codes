module four_to_one(I0,I1,I2,I3,S0,S1,Y);
input I0,I1,I2,I3,S0,S1;
output Y;
wire w1,w2,w3,w4,w5,w6;
not n1(w1,S0);
not n2(w2,S1);
and a1(w3,w1,w2,I0);
and a2(w4,w1,S1,I1);
and a3(w5,S0,w2,I2);
and a4(w6,S0,S1,I3);
or o1(Y,w3,w4,w5,w6);
endmodule
module big_mux(S0,S1,S2,S3,I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,Out);
input S0,S1,S2,S3,I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15;
output Out;
wire q1,q2,q3,q4,q5;
four_to_one f1(I0,I1,I2,I3,S0,S1,q1);
four_to_one f2(I4,I5,I6,I7,S0,S1,q2);
four_to_one f3(I8,I9,I10,I11,S0,S1,q3);
four_to_one f4(I12,I13,I14,I15,S0,S1,q4);
four_to_one f5(q1,q2,q3,q4,S2,S3,Out);
endmodule
module big_mux_tb;
reg S0,S1,S2,S3,I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15;
wire Out;
big_mux b1(S0,S1,S2,S3,I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,Out);
initial
begin
    S0=0;S1=0;S2=0;S3=0;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    $monitor("Time=%0t,S0=%b,S1=%b,S2=%b,S3=%b,I0=%b,I1=%b,I2=%b,I3=%b,I4=%b,I5=%b,I6=%b,I7=%b,I8=%b,I9=%b,I10=%b,I11=%b,I12=%b,I13=%b,I14=%b,I15=%b,Out=%b",$time,S0,S1,S2,S3,I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,Out);
    #10 S0=0;S1=0;S2=0;S3=1;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=0;S1=0;S2=1;S3=0;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=0;S1=0;S2=1;S3=1;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=0;S1=1;S2=0;S3=0;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=0;S1=1;S2=0;S3=1;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=0;S1=1;S2=1;S3=0;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=0;S1=1;S2=1;S3=1;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=1;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=1;S1=0;S2=0;S3=0;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=1;S1=0;S2=0;S3=1;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=1;S1=0;S2=1;S3=0;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=1;S1=0;S2=1;S3=1;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=1;S1=1;S2=0;S3=0;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=1;S1=1;S2=0;S3=1;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=0;I14=0;I15=0;
    #10 S0=1;S1=1;S2=1;S3=0;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
    #10 S0=1;S1=1;S2=1;S3=1;I0=1;I1=0;I2=0;I3=1;I4=0;I5=1;I6=1;I7=0;I8=0;I9=1;I10=0;I11=0;I12=1;I13=1;I14=0;I15=0;
end
endmodule